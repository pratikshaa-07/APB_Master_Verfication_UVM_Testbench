`include "uvm_macros.svh"

package apb_pkg;
import uvm_pkg::*;
//  `include "uvm_pkg.sv"
  //`include "morse_defines.sv"
  `include "seq_item.sv"
  `include "sequence.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "active_monitor.sv"
  `include "passive_monitor.sv"
  `include "active_agent.sv"
  `include "passive_agent.sv"
  `include "scoreboard.sv"
  `include "subscriber.sv"
  `include "environment.sv"
  `include "test.sv"
endpackage

